`timescale 1ns / 1ps

module beer_draft_top(
    clk,
    reset,
    next,draft,
    beer_level,
    beer, 
    state_display);
        
      // WRITE LOGIC HERE
        

endmodule
